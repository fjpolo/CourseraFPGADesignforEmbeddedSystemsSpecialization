-- nios_sys.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_sys is
	port (
		clk_clk                   : in  std_logic                    := '0';             --                clk.clk
		pio_button_export         : in  std_logic                    := '0';             --         pio_button.export
		pio_leds_export           : out std_logic_vector(7 downto 0);                    --           pio_leds.export
		pio_lis3dh_export         : in  std_logic_vector(1 downto 0) := (others => '0'); --         pio_lis3dh.export
		pll_locked_conduit_export : out std_logic;                                       -- pll_locked_conduit.export
		reset_reset_n             : in  std_logic                    := '0';             --              reset.reset_n
		spi_lis3dh_MISO           : in  std_logic                    := '0';             --         spi_lis3dh.MISO
		spi_lis3dh_MOSI           : out std_logic;                                       --                   .MOSI
		spi_lis3dh_SCLK           : out std_logic;                                       --                   .SCLK
		spi_lis3dh_SS_n           : out std_logic                                        --                   .SS_n
	);
end entity nios_sys;

architecture rtl of nios_sys is
	component nios_sys_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_sys_jtag_uart;

	component nios_sys_nios is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(16 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(16 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_sys_nios;

	component nios_sys_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios_sys_onchip_ram;

	component nios_sys_pio_button is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_sys_pio_button;

	component nios_sys_pio_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios_sys_pio_leds;

	component nios_sys_pio_lis3dh is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_sys_pio_lis3dh;

	component nios_sys_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component nios_sys_pll;

	component nios_sys_spi_lis3dh is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component nios_sys_spi_lis3dh;

	component nios_sys_sys_id is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_sys_sys_id;

	component nios_sys_mm_interconnect_0 is
		port (
			clk12mhz_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			nios_reset_reset_bridge_in_reset_reset                : in  std_logic                     := 'X';             -- reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios_data_master_address                              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios_data_master_waitrequest                          : out std_logic;                                        -- waitrequest
			nios_data_master_byteenable                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios_data_master_read                                 : in  std_logic                     := 'X';             -- read
			nios_data_master_readdata                             : out std_logic_vector(31 downto 0);                    -- readdata
			nios_data_master_write                                : in  std_logic                     := 'X';             -- write
			nios_data_master_writedata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios_data_master_debugaccess                          : in  std_logic                     := 'X';             -- debugaccess
			nios_instruction_master_address                       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios_instruction_master_waitrequest                   : out std_logic;                                        -- waitrequest
			nios_instruction_master_read                          : in  std_logic                     := 'X';             -- read
			nios_instruction_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			nios_debug_mem_slave_address                          : out std_logic_vector(8 downto 0);                     -- address
			nios_debug_mem_slave_write                            : out std_logic;                                        -- write
			nios_debug_mem_slave_read                             : out std_logic;                                        -- read
			nios_debug_mem_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_debug_mem_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			nios_debug_mem_slave_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			nios_debug_mem_slave_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			nios_debug_mem_slave_debugaccess                      : out std_logic;                                        -- debugaccess
			onchip_ram_s1_address                                 : out std_logic_vector(12 downto 0);                    -- address
			onchip_ram_s1_write                                   : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                   : out std_logic;                                        -- clken
			pio_button_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_button_s1_write                                   : out std_logic;                                        -- write
			pio_button_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_button_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			pio_button_s1_chipselect                              : out std_logic;                                        -- chipselect
			pio_leds_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			pio_leds_s1_write                                     : out std_logic;                                        -- write
			pio_leds_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_leds_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			pio_leds_s1_chipselect                                : out std_logic;                                        -- chipselect
			pio_lis3dh_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_lis3dh_s1_write                                   : out std_logic;                                        -- write
			pio_lis3dh_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_lis3dh_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			pio_lis3dh_s1_chipselect                              : out std_logic;                                        -- chipselect
			pll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_pll_slave_write                                   : out std_logic;                                        -- write
			pll_pll_slave_read                                    : out std_logic;                                        -- read
			pll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			spi_lis3dh_spi_control_port_address                   : out std_logic_vector(2 downto 0);                     -- address
			spi_lis3dh_spi_control_port_write                     : out std_logic;                                        -- write
			spi_lis3dh_spi_control_port_read                      : out std_logic;                                        -- read
			spi_lis3dh_spi_control_port_readdata                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_lis3dh_spi_control_port_writedata                 : out std_logic_vector(15 downto 0);                    -- writedata
			spi_lis3dh_spi_control_port_chipselect                : out std_logic;                                        -- chipselect
			sys_id_control_slave_address                          : out std_logic_vector(0 downto 0);                     -- address
			sys_id_control_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component nios_sys_mm_interconnect_0;

	component nios_sys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_sys_irq_mapper;

	component nios_sys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_sys_rst_controller;

	component nios_sys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_sys_rst_controller_001;

	signal pll_c0_clk                                                    : std_logic;                     -- pll:c0 -> [irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_c0_clk, nios:clk, onchip_ram:clk, pio_button:clk, pio_leds:clk, pio_lis3dh:clk, rst_controller:clk, spi_lis3dh:clk, sys_id:clock]
	signal nios_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	signal nios_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	signal nios_data_master_debugaccess                                  : std_logic;                     -- nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	signal nios_data_master_address                                      : std_logic_vector(16 downto 0); -- nios:d_address -> mm_interconnect_0:nios_data_master_address
	signal nios_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	signal nios_data_master_read                                         : std_logic;                     -- nios:d_read -> mm_interconnect_0:nios_data_master_read
	signal nios_data_master_write                                        : std_logic;                     -- nios:d_write -> mm_interconnect_0:nios_data_master_write
	signal nios_data_master_writedata                                    : std_logic_vector(31 downto 0); -- nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	signal nios_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	signal nios_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	signal nios_instruction_master_address                               : std_logic_vector(16 downto 0); -- nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	signal nios_instruction_master_read                                  : std_logic;                     -- nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sys_id_control_slave_readdata               : std_logic_vector(31 downto 0); -- sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	signal mm_interconnect_0_sys_id_control_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	signal mm_interconnect_0_nios_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	signal mm_interconnect_0_nios_debug_mem_slave_waitrequest            : std_logic;                     -- nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	signal mm_interconnect_0_nios_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	signal mm_interconnect_0_nios_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	signal mm_interconnect_0_nios_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                      : std_logic_vector(31 downto 0); -- pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_pll_slave_address -> pll:address
	signal mm_interconnect_0_pll_pll_slave_read                          : std_logic;                     -- mm_interconnect_0:pll_pll_slave_read -> pll:read
	signal mm_interconnect_0_pll_pll_slave_write                         : std_logic;                     -- mm_interconnect_0:pll_pll_slave_write -> pll:write
	signal mm_interconnect_0_pll_pll_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	signal mm_interconnect_0_onchip_ram_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                       : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_pio_lis3dh_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:pio_lis3dh_s1_chipselect -> pio_lis3dh:chipselect
	signal mm_interconnect_0_pio_lis3dh_s1_readdata                      : std_logic_vector(31 downto 0); -- pio_lis3dh:readdata -> mm_interconnect_0:pio_lis3dh_s1_readdata
	signal mm_interconnect_0_pio_lis3dh_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_lis3dh_s1_address -> pio_lis3dh:address
	signal mm_interconnect_0_pio_lis3dh_s1_write                         : std_logic;                     -- mm_interconnect_0:pio_lis3dh_s1_write -> mm_interconnect_0_pio_lis3dh_s1_write:in
	signal mm_interconnect_0_pio_lis3dh_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_lis3dh_s1_writedata -> pio_lis3dh:writedata
	signal mm_interconnect_0_pio_leds_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pio_leds_s1_chipselect -> pio_leds:chipselect
	signal mm_interconnect_0_pio_leds_s1_readdata                        : std_logic_vector(31 downto 0); -- pio_leds:readdata -> mm_interconnect_0:pio_leds_s1_readdata
	signal mm_interconnect_0_pio_leds_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_leds_s1_address -> pio_leds:address
	signal mm_interconnect_0_pio_leds_s1_write                           : std_logic;                     -- mm_interconnect_0:pio_leds_s1_write -> mm_interconnect_0_pio_leds_s1_write:in
	signal mm_interconnect_0_pio_leds_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_leds_s1_writedata -> pio_leds:writedata
	signal mm_interconnect_0_pio_button_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:pio_button_s1_chipselect -> pio_button:chipselect
	signal mm_interconnect_0_pio_button_s1_readdata                      : std_logic_vector(31 downto 0); -- pio_button:readdata -> mm_interconnect_0:pio_button_s1_readdata
	signal mm_interconnect_0_pio_button_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_button_s1_address -> pio_button:address
	signal mm_interconnect_0_pio_button_s1_write                         : std_logic;                     -- mm_interconnect_0:pio_button_s1_write -> mm_interconnect_0_pio_button_s1_write:in
	signal mm_interconnect_0_pio_button_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_button_s1_writedata -> pio_button:writedata
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:spi_lis3dh_spi_control_port_chipselect -> spi_lis3dh:spi_select
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_readdata        : std_logic_vector(15 downto 0); -- spi_lis3dh:data_to_cpu -> mm_interconnect_0:spi_lis3dh_spi_control_port_readdata
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_lis3dh_spi_control_port_address -> spi_lis3dh:mem_addr
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_read            : std_logic;                     -- mm_interconnect_0:spi_lis3dh_spi_control_port_read -> mm_interconnect_0_spi_lis3dh_spi_control_port_read:in
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_write           : std_logic;                     -- mm_interconnect_0:spi_lis3dh_spi_control_port_write -> mm_interconnect_0_spi_lis3dh_spi_control_port_write:in
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_writedata       : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_lis3dh_spi_control_port_writedata -> spi_lis3dh:data_from_cpu
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- spi_lis3dh:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- pio_lis3dh:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- pio_button:irq -> irq_mapper:receiver3_irq
	signal nios_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [nios:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	signal nios_debug_reset_request_reset                                : std_logic;                     -- nios:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_pio_lis3dh_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_pio_lis3dh_s1_write:inv -> pio_lis3dh:write_n
	signal mm_interconnect_0_pio_leds_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_leds_s1_write:inv -> pio_leds:write_n
	signal mm_interconnect_0_pio_button_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_pio_button_s1_write:inv -> pio_button:write_n
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_spi_lis3dh_spi_control_port_read:inv -> spi_lis3dh:read_n
	signal mm_interconnect_0_spi_lis3dh_spi_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_spi_lis3dh_spi_control_port_write:inv -> spi_lis3dh:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart:rst_n, nios:reset_n, pio_button:reset_n, pio_leds:reset_n, pio_lis3dh:reset_n, spi_lis3dh:reset_n, sys_id:reset_n]

begin

	jtag_uart : component nios_sys_jtag_uart
		port map (
			clk            => pll_c0_clk,                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	nios : component nios_sys_nios
		port map (
			clk                                 => pll_c0_clk,                                         --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,           --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                 --                          .reset_req
			d_address                           => nios_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_data_master_read,                              --                          .read
			d_readdata                          => nios_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_data_master_write,                             --                          .write
			d_writedata                         => nios_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_instruction_master_read,                       --                          .read
			i_readdata                          => nios_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                -- custom_instruction_master.readra
		);

	onchip_ram : component nios_sys_onchip_ram
		port map (
			clk        => pll_c0_clk,                                 --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pio_button : component nios_sys_pio_button
		port map (
			clk        => pll_c0_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_pio_button_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_button_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_button_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_button_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_button_s1_readdata,        --                    .readdata
			in_port    => pio_button_export,                               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                         --                 irq.irq
		);

	pio_leds : component nios_sys_pio_leds
		port map (
			clk        => pll_c0_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_leds_s1_readdata,        --                    .readdata
			out_port   => pio_leds_export                                -- external_connection.export
		);

	pio_lis3dh : component nios_sys_pio_lis3dh
		port map (
			clk        => pll_c0_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_pio_lis3dh_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_lis3dh_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_lis3dh_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_lis3dh_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_lis3dh_s1_readdata,        --                    .readdata
			in_port    => pio_lis3dh_export,                               -- external_connection.export
			irq        => irq_mapper_receiver2_irq                         --                 irq.irq
		);

	pll : component nios_sys_pll
		port map (
			clk                => clk_clk,                                   --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			locked             => pll_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			c1                 => open,                                      --           (terminated)
			c2                 => open,                                      --           (terminated)
			c3                 => open,                                      --           (terminated)
			c4                 => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "000",                                     --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	spi_lis3dh : component nios_sys_spi_lis3dh
		port map (
			clk           => pll_c0_clk,                                                    --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                      --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_lis3dh_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_lis3dh_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_lis3dh_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_lis3dh_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_lis3dh_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_lis3dh_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver0_irq,                                      --              irq.irq
			MISO          => spi_lis3dh_MISO,                                               --         external.export
			MOSI          => spi_lis3dh_MOSI,                                               --                 .export
			SCLK          => spi_lis3dh_SCLK,                                               --                 .export
			SS_n          => spi_lis3dh_SS_n                                                --                 .export
		);

	sys_id : component nios_sys_sys_id
		port map (
			clock    => pll_c0_clk,                                        --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_0_sys_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sys_id_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component nios_sys_mm_interconnect_0
		port map (
			clk12mhz_clk_clk                                      => clk_clk,                                                   --                                    clk12mhz_clk.clk
			pll_c0_clk                                            => pll_c0_clk,                                                --                                          pll_c0.clk
			nios_reset_reset_bridge_in_reset_reset                => rst_controller_reset_out_reset,                            --                nios_reset_reset_bridge_in_reset.reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                        -- pll_inclk_interface_reset_reset_bridge_in_reset.reset
			nios_data_master_address                              => nios_data_master_address,                                  --                                nios_data_master.address
			nios_data_master_waitrequest                          => nios_data_master_waitrequest,                              --                                                .waitrequest
			nios_data_master_byteenable                           => nios_data_master_byteenable,                               --                                                .byteenable
			nios_data_master_read                                 => nios_data_master_read,                                     --                                                .read
			nios_data_master_readdata                             => nios_data_master_readdata,                                 --                                                .readdata
			nios_data_master_write                                => nios_data_master_write,                                    --                                                .write
			nios_data_master_writedata                            => nios_data_master_writedata,                                --                                                .writedata
			nios_data_master_debugaccess                          => nios_data_master_debugaccess,                              --                                                .debugaccess
			nios_instruction_master_address                       => nios_instruction_master_address,                           --                         nios_instruction_master.address
			nios_instruction_master_waitrequest                   => nios_instruction_master_waitrequest,                       --                                                .waitrequest
			nios_instruction_master_read                          => nios_instruction_master_read,                              --                                                .read
			nios_instruction_master_readdata                      => nios_instruction_master_readdata,                          --                                                .readdata
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                                .chipselect
			nios_debug_mem_slave_address                          => mm_interconnect_0_nios_debug_mem_slave_address,            --                            nios_debug_mem_slave.address
			nios_debug_mem_slave_write                            => mm_interconnect_0_nios_debug_mem_slave_write,              --                                                .write
			nios_debug_mem_slave_read                             => mm_interconnect_0_nios_debug_mem_slave_read,               --                                                .read
			nios_debug_mem_slave_readdata                         => mm_interconnect_0_nios_debug_mem_slave_readdata,           --                                                .readdata
			nios_debug_mem_slave_writedata                        => mm_interconnect_0_nios_debug_mem_slave_writedata,          --                                                .writedata
			nios_debug_mem_slave_byteenable                       => mm_interconnect_0_nios_debug_mem_slave_byteenable,         --                                                .byteenable
			nios_debug_mem_slave_waitrequest                      => mm_interconnect_0_nios_debug_mem_slave_waitrequest,        --                                                .waitrequest
			nios_debug_mem_slave_debugaccess                      => mm_interconnect_0_nios_debug_mem_slave_debugaccess,        --                                                .debugaccess
			onchip_ram_s1_address                                 => mm_interconnect_0_onchip_ram_s1_address,                   --                                   onchip_ram_s1.address
			onchip_ram_s1_write                                   => mm_interconnect_0_onchip_ram_s1_write,                     --                                                .write
			onchip_ram_s1_readdata                                => mm_interconnect_0_onchip_ram_s1_readdata,                  --                                                .readdata
			onchip_ram_s1_writedata                               => mm_interconnect_0_onchip_ram_s1_writedata,                 --                                                .writedata
			onchip_ram_s1_byteenable                              => mm_interconnect_0_onchip_ram_s1_byteenable,                --                                                .byteenable
			onchip_ram_s1_chipselect                              => mm_interconnect_0_onchip_ram_s1_chipselect,                --                                                .chipselect
			onchip_ram_s1_clken                                   => mm_interconnect_0_onchip_ram_s1_clken,                     --                                                .clken
			pio_button_s1_address                                 => mm_interconnect_0_pio_button_s1_address,                   --                                   pio_button_s1.address
			pio_button_s1_write                                   => mm_interconnect_0_pio_button_s1_write,                     --                                                .write
			pio_button_s1_readdata                                => mm_interconnect_0_pio_button_s1_readdata,                  --                                                .readdata
			pio_button_s1_writedata                               => mm_interconnect_0_pio_button_s1_writedata,                 --                                                .writedata
			pio_button_s1_chipselect                              => mm_interconnect_0_pio_button_s1_chipselect,                --                                                .chipselect
			pio_leds_s1_address                                   => mm_interconnect_0_pio_leds_s1_address,                     --                                     pio_leds_s1.address
			pio_leds_s1_write                                     => mm_interconnect_0_pio_leds_s1_write,                       --                                                .write
			pio_leds_s1_readdata                                  => mm_interconnect_0_pio_leds_s1_readdata,                    --                                                .readdata
			pio_leds_s1_writedata                                 => mm_interconnect_0_pio_leds_s1_writedata,                   --                                                .writedata
			pio_leds_s1_chipselect                                => mm_interconnect_0_pio_leds_s1_chipselect,                  --                                                .chipselect
			pio_lis3dh_s1_address                                 => mm_interconnect_0_pio_lis3dh_s1_address,                   --                                   pio_lis3dh_s1.address
			pio_lis3dh_s1_write                                   => mm_interconnect_0_pio_lis3dh_s1_write,                     --                                                .write
			pio_lis3dh_s1_readdata                                => mm_interconnect_0_pio_lis3dh_s1_readdata,                  --                                                .readdata
			pio_lis3dh_s1_writedata                               => mm_interconnect_0_pio_lis3dh_s1_writedata,                 --                                                .writedata
			pio_lis3dh_s1_chipselect                              => mm_interconnect_0_pio_lis3dh_s1_chipselect,                --                                                .chipselect
			pll_pll_slave_address                                 => mm_interconnect_0_pll_pll_slave_address,                   --                                   pll_pll_slave.address
			pll_pll_slave_write                                   => mm_interconnect_0_pll_pll_slave_write,                     --                                                .write
			pll_pll_slave_read                                    => mm_interconnect_0_pll_pll_slave_read,                      --                                                .read
			pll_pll_slave_readdata                                => mm_interconnect_0_pll_pll_slave_readdata,                  --                                                .readdata
			pll_pll_slave_writedata                               => mm_interconnect_0_pll_pll_slave_writedata,                 --                                                .writedata
			spi_lis3dh_spi_control_port_address                   => mm_interconnect_0_spi_lis3dh_spi_control_port_address,     --                     spi_lis3dh_spi_control_port.address
			spi_lis3dh_spi_control_port_write                     => mm_interconnect_0_spi_lis3dh_spi_control_port_write,       --                                                .write
			spi_lis3dh_spi_control_port_read                      => mm_interconnect_0_spi_lis3dh_spi_control_port_read,        --                                                .read
			spi_lis3dh_spi_control_port_readdata                  => mm_interconnect_0_spi_lis3dh_spi_control_port_readdata,    --                                                .readdata
			spi_lis3dh_spi_control_port_writedata                 => mm_interconnect_0_spi_lis3dh_spi_control_port_writedata,   --                                                .writedata
			spi_lis3dh_spi_control_port_chipselect                => mm_interconnect_0_spi_lis3dh_spi_control_port_chipselect,  --                                                .chipselect
			sys_id_control_slave_address                          => mm_interconnect_0_sys_id_control_slave_address,            --                            sys_id_control_slave.address
			sys_id_control_slave_readdata                         => mm_interconnect_0_sys_id_control_slave_readdata            --                                                .readdata
		);

	irq_mapper : component nios_sys_irq_mapper
		port map (
			clk           => pll_c0_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios_irq_irq                    --    sender.irq
		);

	rst_controller : component nios_sys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios_debug_reset_request_reset,     -- reset_in1.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component nios_sys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios_debug_reset_request_reset,     -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_pio_lis3dh_s1_write_ports_inv <= not mm_interconnect_0_pio_lis3dh_s1_write;

	mm_interconnect_0_pio_leds_s1_write_ports_inv <= not mm_interconnect_0_pio_leds_s1_write;

	mm_interconnect_0_pio_button_s1_write_ports_inv <= not mm_interconnect_0_pio_button_s1_write;

	mm_interconnect_0_spi_lis3dh_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_lis3dh_spi_control_port_read;

	mm_interconnect_0_spi_lis3dh_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_lis3dh_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_sys
